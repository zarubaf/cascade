/*
Copyright 2010, D. E. Shaw Research.
All rights reserved.

Redistribution and use in source and binary forms, with or without
modification, are permitted provided that the following conditions are
met:

* Redistributions of source code must retain the above copyright
  notice, this list of conditions, and the following disclaimer.

* Redistributions in binary form must reproduce the above copyright
  notice, this list of conditions, and the following disclaimer in the
  documentation and/or other materials provided with the distribution.

* Neither the name of D. E. Shaw Research nor the names of its
  contributors may be used to endorse or promote products derived from
  this software without specific prior written permission.

THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS
"AS IS" AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT
LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR
A PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT
OWNER OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL,
SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT
LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES; LOSS OF USE,
DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY
THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
(INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE
OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
*/

/////////////////////////////////////////////////////////////////
//
// dpi.svh
//
// Copyright (C) 2010 D. E. Shaw Research
//
// Author:  J.P. Grossman (jp.grossman@deshawresearch.com)
// Created: 2/18/2010
//
// `include this file from Verilog in order to use the DPI
// functions.
//
/////////////////////////////////////////////////////////////////

//
// setCModuleParam()
//
// Call this function zero or more times before createCModule to
// set the values of the CModule parameters.
//
import "DPI-C" function void setCModuleParam (input string name, input int value);

//
// createCModule()
//
// Call this function within a wrapper module in order to instantiate
// a CModule and bind its ports to the wrapper's ports.  Sample usage:
//
//     module cmodule_wrapper (<ports>);
//
//         chandle cmodule;
//         initial begin
//             string s;
//             $sformat(s, "%m");
//             cmodule = createCModule("adder", s);
//         end
//
//         <PUSH/POP macros>
//
//     endmodule
//
//
import "DPI-C" function chandle createCModule (input string name, input string verilogName);

//
// clockCModule()
//
// Don't call this function directly; use the `CLOCK_CMODULE macro after the `PUSH_TO_C
// macros and before the `POP_FROM_C macros (Currently the `CLOCK_CMODULE macro just
// calls clockCModule(), but at some point it might perform additional tasks).
//
import "DPI-C" function void clockCModule (input chandle scope, input string clockName);
`define CLOCK_CMODULE(clockName) clockCModule(cmodule, "clockName");

//
// setCModuleTraces()
//
// Enables tracing within the CModules.  Takes a single string argument,
// which is a semicolon-delimited list of trace speciers.  Refer to the
// Cascade documentation for the format of the trace specifiers.
//
import "DPI-C" function void setCModuleTraces (input string traces);

//
// dumpCModuleVars()
//
// Create waves from the Cmodule signals.  Takes a single string argument,
// which is a semicolon-delimited list of dump speciers.  Refer to the
// Cascade documentation for the format of the dump specifiers.
// This must be called before the simulation begins.
//
import "DPI-C" function void dumpCModuleVars (input string dumps);

//
// disableCAssertion()
//
// Disable an assertion within the CModules.  If 'message' matches any substring
// of the error output, then the assertion is ignored.  'message' can contain the
// * and ? wildcards (so $disable_assertion("*") disables all assertions).
//
import "DPI-C" function void disableCAssertion (input string message);

//
// setCParameter()
//
// Set one of the C++ parameters to the specified value.
//
import "DPI-C" function void setCParameter (input string name, input string value);

//
// Functions and macros used to skip over ports when using multiple clocks
//
import "DPI-C" function void ignoreCPort (input chandle scope, input string name, input int isInput);
`define IGNORE_TO_C(port)   ignoreCPort(cmodule, "port", 1);
`define IGNORE_FROM_C(port) ignoreCPort(cmodule, "port", 0);

/***** Functions + Macros Generated by the following program *****

#include <stdio.h>

int main (void)
{
    int i;

    for (i = 32 ; i <= 1024 ; i += 32)
        printf("import \"DPI-C\" function void pushToC%-3d (input chandle scope, input bit [%d:0] b, input string portName, input int sizeInBits);\n", i, i-1);

    printf("\n");
    for (i = 32 ; i <= 1024 ; i += 32)
        printf("import \"DPI-C\" function void popFromC%-3d (input chandle scope, output bit [%d:0] b, input string portName, input int sizeInBits);\n", i, i-1);

    printf("\n`define PUSH_TO_C(port) \\\n");
    printf("if      ($bits(port) <= 32 ) pushToC32 (cmodule, port, \"port\", $bits(port)); \\\n");
    for (i = 64 ; i < 1024 ; i += 32)
        printf("else if ($bits(port) <= %-3d) pushToC%-3d(cmodule, port, \"port\", $bits(port)); \\\n", i, i);
    printf("else                        pushToC1024(cmodule, port, \"port\", $bits(port))\n");

    printf("\n`define POP_FROM_C(port) \\\n");
    printf("begin \\\n");
    printf("    logic [$bits(port)-1:0] tmp_``port; \\\n");
    printf("    if      ($bits(port) <= 32 ) popFromC32 (cmodule, tmp_``port, \"port\", $bits(port)); \\\n");
    for (i = 64 ; i < 1024 ; i += 32)
        printf("    else if ($bits(port) <= %-3d) popFromC%-3d(cmodule, tmp_``port, \"port\", $bits(port)); \\\n", i, i);
    printf("    else                         popFromC1024(cmodule, tmp_``port, \"port\", $bits(port)); \\\n");
    printf("    port <= tmp_``port; \\\n");
    printf("end\n");
}

*****************************************************************/

import "DPI-C" function void pushToC32  (input chandle scope, input bit [31:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void pushToC64  (input chandle scope, input bit [63:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void pushToC96  (input chandle scope, input bit [95:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void pushToC128 (input chandle scope, input bit [127:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void pushToC160 (input chandle scope, input bit [159:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void pushToC192 (input chandle scope, input bit [191:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void pushToC224 (input chandle scope, input bit [223:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void pushToC256 (input chandle scope, input bit [255:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void pushToC288 (input chandle scope, input bit [287:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void pushToC320 (input chandle scope, input bit [319:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void pushToC352 (input chandle scope, input bit [351:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void pushToC384 (input chandle scope, input bit [383:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void pushToC416 (input chandle scope, input bit [415:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void pushToC448 (input chandle scope, input bit [447:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void pushToC480 (input chandle scope, input bit [479:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void pushToC512 (input chandle scope, input bit [511:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void pushToC544 (input chandle scope, input bit [543:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void pushToC576 (input chandle scope, input bit [575:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void pushToC608 (input chandle scope, input bit [607:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void pushToC640 (input chandle scope, input bit [639:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void pushToC672 (input chandle scope, input bit [671:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void pushToC704 (input chandle scope, input bit [703:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void pushToC736 (input chandle scope, input bit [735:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void pushToC768 (input chandle scope, input bit [767:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void pushToC800 (input chandle scope, input bit [799:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void pushToC832 (input chandle scope, input bit [831:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void pushToC864 (input chandle scope, input bit [863:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void pushToC896 (input chandle scope, input bit [895:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void pushToC928 (input chandle scope, input bit [927:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void pushToC960 (input chandle scope, input bit [959:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void pushToC992 (input chandle scope, input bit [991:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void pushToC1024 (input chandle scope, input bit [1023:0] b, input string portName, input int sizeInBits);

import "DPI-C" function void popFromC32  (input chandle scope, output bit [31:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void popFromC64  (input chandle scope, output bit [63:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void popFromC96  (input chandle scope, output bit [95:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void popFromC128 (input chandle scope, output bit [127:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void popFromC160 (input chandle scope, output bit [159:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void popFromC192 (input chandle scope, output bit [191:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void popFromC224 (input chandle scope, output bit [223:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void popFromC256 (input chandle scope, output bit [255:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void popFromC288 (input chandle scope, output bit [287:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void popFromC320 (input chandle scope, output bit [319:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void popFromC352 (input chandle scope, output bit [351:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void popFromC384 (input chandle scope, output bit [383:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void popFromC416 (input chandle scope, output bit [415:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void popFromC448 (input chandle scope, output bit [447:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void popFromC480 (input chandle scope, output bit [479:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void popFromC512 (input chandle scope, output bit [511:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void popFromC544 (input chandle scope, output bit [543:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void popFromC576 (input chandle scope, output bit [575:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void popFromC608 (input chandle scope, output bit [607:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void popFromC640 (input chandle scope, output bit [639:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void popFromC672 (input chandle scope, output bit [671:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void popFromC704 (input chandle scope, output bit [703:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void popFromC736 (input chandle scope, output bit [735:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void popFromC768 (input chandle scope, output bit [767:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void popFromC800 (input chandle scope, output bit [799:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void popFromC832 (input chandle scope, output bit [831:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void popFromC864 (input chandle scope, output bit [863:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void popFromC896 (input chandle scope, output bit [895:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void popFromC928 (input chandle scope, output bit [927:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void popFromC960 (input chandle scope, output bit [959:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void popFromC992 (input chandle scope, output bit [991:0] b, input string portName, input int sizeInBits);
import "DPI-C" function void popFromC1024 (input chandle scope, output bit [1023:0] b, input string portName, input int sizeInBits);

`define PUSH_TO_C(port) \
if      ($bits(port) <= 32 ) pushToC32 (cmodule, port, "port", $bits(port)); \
else if ($bits(port) <= 64 ) pushToC64 (cmodule, port, "port", $bits(port)); \
else if ($bits(port) <= 96 ) pushToC96 (cmodule, port, "port", $bits(port)); \
else if ($bits(port) <= 128) pushToC128(cmodule, port, "port", $bits(port)); \
else if ($bits(port) <= 160) pushToC160(cmodule, port, "port", $bits(port)); \
else if ($bits(port) <= 192) pushToC192(cmodule, port, "port", $bits(port)); \
else if ($bits(port) <= 224) pushToC224(cmodule, port, "port", $bits(port)); \
else if ($bits(port) <= 256) pushToC256(cmodule, port, "port", $bits(port)); \
else if ($bits(port) <= 288) pushToC288(cmodule, port, "port", $bits(port)); \
else if ($bits(port) <= 320) pushToC320(cmodule, port, "port", $bits(port)); \
else if ($bits(port) <= 352) pushToC352(cmodule, port, "port", $bits(port)); \
else if ($bits(port) <= 384) pushToC384(cmodule, port, "port", $bits(port)); \
else if ($bits(port) <= 416) pushToC416(cmodule, port, "port", $bits(port)); \
else if ($bits(port) <= 448) pushToC448(cmodule, port, "port", $bits(port)); \
else if ($bits(port) <= 480) pushToC480(cmodule, port, "port", $bits(port)); \
else if ($bits(port) <= 512) pushToC512(cmodule, port, "port", $bits(port)); \
else if ($bits(port) <= 544) pushToC544(cmodule, port, "port", $bits(port)); \
else if ($bits(port) <= 576) pushToC576(cmodule, port, "port", $bits(port)); \
else if ($bits(port) <= 608) pushToC608(cmodule, port, "port", $bits(port)); \
else if ($bits(port) <= 640) pushToC640(cmodule, port, "port", $bits(port)); \
else if ($bits(port) <= 672) pushToC672(cmodule, port, "port", $bits(port)); \
else if ($bits(port) <= 704) pushToC704(cmodule, port, "port", $bits(port)); \
else if ($bits(port) <= 736) pushToC736(cmodule, port, "port", $bits(port)); \
else if ($bits(port) <= 768) pushToC768(cmodule, port, "port", $bits(port)); \
else if ($bits(port) <= 800) pushToC800(cmodule, port, "port", $bits(port)); \
else if ($bits(port) <= 832) pushToC832(cmodule, port, "port", $bits(port)); \
else if ($bits(port) <= 864) pushToC864(cmodule, port, "port", $bits(port)); \
else if ($bits(port) <= 896) pushToC896(cmodule, port, "port", $bits(port)); \
else if ($bits(port) <= 928) pushToC928(cmodule, port, "port", $bits(port)); \
else if ($bits(port) <= 960) pushToC960(cmodule, port, "port", $bits(port)); \
else if ($bits(port) <= 992) pushToC992(cmodule, port, "port", $bits(port)); \
else                        pushToC1024(cmodule, port, "port", $bits(port));

`define POP_FROM_C(port) \
begin \
    logic [$bits(port)-1:0] tmp_``port; \
    if      ($bits(port) <= 32 ) popFromC32 (cmodule, tmp_``port, "port", $bits(port)); \
    else if ($bits(port) <= 64 ) popFromC64 (cmodule, tmp_``port, "port", $bits(port)); \
    else if ($bits(port) <= 96 ) popFromC96 (cmodule, tmp_``port, "port", $bits(port)); \
    else if ($bits(port) <= 128) popFromC128(cmodule, tmp_``port, "port", $bits(port)); \
    else if ($bits(port) <= 160) popFromC160(cmodule, tmp_``port, "port", $bits(port)); \
    else if ($bits(port) <= 192) popFromC192(cmodule, tmp_``port, "port", $bits(port)); \
    else if ($bits(port) <= 224) popFromC224(cmodule, tmp_``port, "port", $bits(port)); \
    else if ($bits(port) <= 256) popFromC256(cmodule, tmp_``port, "port", $bits(port)); \
    else if ($bits(port) <= 288) popFromC288(cmodule, tmp_``port, "port", $bits(port)); \
    else if ($bits(port) <= 320) popFromC320(cmodule, tmp_``port, "port", $bits(port)); \
    else if ($bits(port) <= 352) popFromC352(cmodule, tmp_``port, "port", $bits(port)); \
    else if ($bits(port) <= 384) popFromC384(cmodule, tmp_``port, "port", $bits(port)); \
    else if ($bits(port) <= 416) popFromC416(cmodule, tmp_``port, "port", $bits(port)); \
    else if ($bits(port) <= 448) popFromC448(cmodule, tmp_``port, "port", $bits(port)); \
    else if ($bits(port) <= 480) popFromC480(cmodule, tmp_``port, "port", $bits(port)); \
    else if ($bits(port) <= 512) popFromC512(cmodule, tmp_``port, "port", $bits(port)); \
    else if ($bits(port) <= 544) popFromC544(cmodule, tmp_``port, "port", $bits(port)); \
    else if ($bits(port) <= 576) popFromC576(cmodule, tmp_``port, "port", $bits(port)); \
    else if ($bits(port) <= 608) popFromC608(cmodule, tmp_``port, "port", $bits(port)); \
    else if ($bits(port) <= 640) popFromC640(cmodule, tmp_``port, "port", $bits(port)); \
    else if ($bits(port) <= 672) popFromC672(cmodule, tmp_``port, "port", $bits(port)); \
    else if ($bits(port) <= 704) popFromC704(cmodule, tmp_``port, "port", $bits(port)); \
    else if ($bits(port) <= 736) popFromC736(cmodule, tmp_``port, "port", $bits(port)); \
    else if ($bits(port) <= 768) popFromC768(cmodule, tmp_``port, "port", $bits(port)); \
    else if ($bits(port) <= 800) popFromC800(cmodule, tmp_``port, "port", $bits(port)); \
    else if ($bits(port) <= 832) popFromC832(cmodule, tmp_``port, "port", $bits(port)); \
    else if ($bits(port) <= 864) popFromC864(cmodule, tmp_``port, "port", $bits(port)); \
    else if ($bits(port) <= 896) popFromC896(cmodule, tmp_``port, "port", $bits(port)); \
    else if ($bits(port) <= 928) popFromC928(cmodule, tmp_``port, "port", $bits(port)); \
    else if ($bits(port) <= 960) popFromC960(cmodule, tmp_``port, "port", $bits(port)); \
    else if ($bits(port) <= 992) popFromC992(cmodule, tmp_``port, "port", $bits(port)); \
    else                         popFromC1024(cmodule, tmp_``port, "port", $bits(port)); \
    port <= tmp_``port; \
end

